/*
 * Copyright (C) 2020 CESNET z. s. p. o.
 * SPDX-License-Identifier: BSD-3-Clause
*/

`include "interface.sv"

package avst_tx;
    `include "config.sv"
    `include "transaction.sv"
    `include "driver.sv"
    `include "agent.sv"
endpackage

/*
 * packet_generator_pkg.sv: SystemVerilog Packet generator package
 * Copyright (C) 2008 CESNET
 * Author(s):  Vlastimil Kosar <xkosar02@stud.fit.vutbr.cz>
 *
 * SPDX-License-Identifier: BSD-3-Clause
 *
 *
 * TODO:
 */

package packet_generator_pkg;
  `include "layer.sv"
  `include "ethernet_II.sv"
  `include "ethernet_II_dotq.sv"
  `include "ethernet_II_dotad.sv"
  `include "icmp.sv"
  `include "icmpv6.sv"
  `include "ipv4.sv"
  `include "ipv6.sv"
  `include "raw.sv"
  `include "raw_pattern.sv"
  `include "tcp.sv"
  `include "udp.sv"
  `include "mpls.sv"
  `include "packetTransaction.sv"
  `include "packetGenerator.sv"
endpackage : packet_generator_pkg

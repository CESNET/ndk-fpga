
/*
 * file       : pkg.sv
 * Copyright (C) 2023 CESNET z. s. p. o.
 * description: probe package
 * date       : 2023
 * author     : Radek Iša <isa@cesnet.ch>
 *
 * SPDX-License-Identifier: BSD-3-Clause
*/

package uvm_probe;

    `include "uvm_macros.svh"
    import uvm_pkg::*;

    `include "data.sv"
    `include "cbs.sv"
    `include "pool.sv"


endpackage

// pkg.sv: Package for pcie
// Copyright (C) 2024 CESNET z. s. p. o.
// Author:  Radek Iša <isa@cesnet.cz>

// SPDX-License-Identifier: BSD-3-Clause

`ifndef PCIE_EXTEND_ENV_SV
`define PCIE_EXTEND_ENV_SV

package uvm_pcie_extend;

    `include "uvm_macros.svh"
    import uvm_pkg::*;

    `include "header.sv"

endpackage

`endif

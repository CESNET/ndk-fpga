//-- tbench.sv: Testbench
//-- Copyright (C) 2022 CESNET z. s. p. o.
//-- Author:   Daniel Kříž <xkrizd01@vutbr.cz>

//-- SPDX-License-Identifier: BSD-3-Clause

import uvm_pkg::*;
`include "uvm_macros.svh"
import test::*;

module testbench;

    // -------------------------------------------------------------------------------------------------------------------------------------------------------------------
    // Signals
    logic CLK = 0;
    logic RST = 0;

    // -------------------------------------------------------------------------------------------------------------------------------------------------------------------
    // Interfaces
    reset_if  reset(CLK);
    mvb_if #(MVB_ITEMS, REG_DEPTH-SLICE_WIDTH) mvb_rx(CLK);
    mvb_if #(MVB_ITEMS, LUT_WIDTH) mvb_tx(CLK);
    mi_if #(SW_WIDTH, REG_DEPTH) mi_config(CLK);

    // -------------------------------------------------------------------------------------------------------------------------------------------------------------------
    // Define clock period
    always #(CLK_PERIOD) CLK = ~CLK;

    // -------------------------------------------------------------------------------------------------------------------------------------------------------------------
    // Initial reset
    initial begin
        RST = 1;
        #(RESET_CLKS*CLK_PERIOD)
        RST = 0;
    end


    // -------------------------------------------------------------------------------------------------------------------------------------------------------------------
    // Start of tests
    initial begin
        uvm_root m_root;
        // Configuration of database
        uvm_config_db#(virtual reset_if)::set(null, "", "vif_reset", reset);
        uvm_config_db#(virtual mvb_if #(MVB_ITEMS, REG_DEPTH-SLICE_WIDTH))::set(null, "", "vif_rx", mvb_rx);
        uvm_config_db#(virtual mvb_if #(MVB_ITEMS, LUT_WIDTH))::set(null, "", "vif_tx", mvb_tx);
        uvm_config_db#(virtual mi_if #(SW_WIDTH, REG_DEPTH))::set(null, "", "vif_mi", mi_config);

        m_root = uvm_root::get();
        m_root.finish_on_completion = 0;
        m_root.set_report_id_action_hier("ILLEGALNAME",UVM_NO_ACTION);

        uvm_config_db#(int)            ::set(null, "", "recording_detail", 0);
        uvm_config_db#(uvm_bitstream_t)::set(null, "", "recording_detail", 0);

        run_test();
        $stop(2);
    end

    // -------------------------------------------------------------------------------------------------------------------------------------------------------------------
    // DUT
    DUT DUT_U (
        .CLK    (CLK),
        .RST    (reset.RESET),
        .mvb_rx (mvb_rx),
        .mvb_tx (mvb_tx),
        .config_mi  (mi_config)
    );

    // -------------------------------------------------------------------------------------------------------------------------------------------------------------------
    // Properties
    // mvb_property #(
    //     .MVB_ITEMS       (MVB_ITEMS),
    //     .ITEM_WIDTH  (ITEM_WIDTH)
    // )
    // property_rd(
    //     .RESET (reset.RESET),
    //     .vif   (mvb_tx)
    // );

    // mvb_property  #(
    //     .MVB_ITEMS      (MVB_ITEMS),
    //     .ITEM_WIDTH (ITEM_WIDTH)
    // )
    // property_wr (
    //     .RESET (reset.RESET),
    //     .vif   (mvb_rx)
    // );

endmodule

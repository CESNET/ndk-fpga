-- This file is only for verification purposes only

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

package combo_user_const is
    constant PCIE_CORE_DEBUG_ENABLE : boolean := false;
    constant PCIE_CTRL_DEBUG_ENABLE : boolean := false;
end combo_user_const;

package body combo_user_const is
end combo_user_const;

/*
 * Copyright (C) 2020 CESNET z. s. p. o.
 * SPDX-License-Identifier: BSD-3-Clause
*/

///////////////////////////////////////////////////////////////////////////////
// configuration file for avalon TX UVM agent
class config_item;

   // Variables
   int unsigned wait_delay = 3;

   // functions
endclass


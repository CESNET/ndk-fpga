
//let min(a,b) = (a < b) ? a : b;

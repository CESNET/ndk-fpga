-- h3_pack.vhd: Package containing available H3 core configurations
-- Copyright (C) 2024 CESNET z. s. p. o.
-- Author(s): Oliver Gurka <oliver.gurka@cesnet.cz>
--
-- SPDX-License-Identifier: BSD-3-Clause

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

package h3_pack is

    type h3_config is record
        tag         : string;
        key_width   : natural;
        hash_width  : natural;
        matrix      : std_logic_vector;
    end record;

    constant H3C_64x16 : h3_config(matrix(64 * 16 - 1 downto 0)) := (
        tag         => "H3C_64x16",
        key_width   => 64,
        hash_width  => 16,
        matrix      => "1111110111101110110101111011011011110101010101111110100001110101001011000110111010101010101101010011110011000011111010001100011011101001011001111111100010000111000110101000110100101001000000100111100001010100111111101101000100000100001101101011011101110000101011111110100001110100111000001010010000011010101000100101101010001110111100100101000010101111010110100000011001100111111111100100011100110111110001110001101010000000001001000111011110111111100000000011011011100000111111011100000110111101110110111010110010101010000011001010101010101001010010011000001111111011010000001000101001000110011001111011001111011100100001010111010010110000110010001001110111001011001111111111101110010100011101000000000110001000000001111110110110000111101111111010011000110110111111011101010001110110001010101111010110001100010010110110001000001101100101000110111010100111001101110010110101100001010001001001101010011010001111010100001101101100110111000111111001101001101010011010011001111000000000001010011000001001110101010011101100101100"
    );

    constant H3C_64x22 : h3_config(matrix(64 * 22 - 1 downto 0)) := (
        tag         => "H3C_64x22",
        key_width   => 64,
        hash_width  => 22,
        matrix      => "1010011101010011010001000011100011101001011010101001010010000100011110000101111011010111000011000101100111000111101001001000100010000110100100010110000010111011101101001101111100110100100001110000001001000010110011010011101000001111111000010000100000100010001001111101101111000000101110101001101011111100010011100010100000010111101010011000011110110011010110111011110111011100000011101011011001101010000100000101011100010000101101010001011100111101111001101110101011111111010001000000010101110101000011001011010100100000101101010100011111001100111101010011000111111010100111101001001111011110101100100000000001011110011101110001010001101000001101111011110000000001101011111111100000010010011110100010101100110010000000010111011101011111010110100010001100001010000110000100010001111100110110101101110000011011101101000110011111100100100111010110101011111111001011101010101101100001101000100101011110101011110110001011000011010011001011000001111110100001110011001001101011011001110111000011110111000101100010001100100000001110001010001001010101100010001110111011010001100111010111110110111011110100010100111010110010011111001100110101111010011011101111011010010110101101101010001000000100101000111011101010101100011111000100010011000001111111001010010100010000110101010110100101010001111011101101110101000010000001000001001001001001110111101101011111110010011011000101110000000101001010110000010001011100101101"
    );

    constant H3C_22x11 : h3_config(matrix(22 * 11 - 1 downto 0)) := (
        tag         => "H3C_22x11",
        key_width   => 22,
        hash_width  => 11,
        matrix      =>"11000000000111101110001100011000001111010111000100010110000010101100101101000000100010101000010001010000110011001101101101010000001110001000010001110100101001111001111100000000110010010000000111000001101010000001000100000011110001101000011010"
    );

    constant H3C_256x64 : h3_config(matrix(256 * 64 - 1 downto 0)) := (
        tag         => "H3C_256x64",
        key_width   => 256,
        hash_width  => 64,
        matrix      => "1111101000101111100100010010010100001110110110100101111101110101100010101100101010001001010111011011010011010100010101101001111111001010011100000011001101010011011000011010101000011011000111100101000101010000101011010010110000110000010011110111010000000110001000000010000100011100101110001110010100100001110011010000100101011001111100110000100001000101111011101011111011100000101010110001010001010010111111011100100001001100011000000110111101001110010010000010100111000001011001101010111011010101001111000111001001101011010110011001001110100110000101101111000100110111100101111111000010001000010001010000011101000100010110110111101111001001100001100010101111011000010011111010001100111000001010000000011001110110100100100101100010110111001111110101101101100111011110101101101010111110010010001011111111000000111011110001011001001011010010101110000111111110010101000101101100110011001110000001011111101010111111010111101110010000100110001110101100110010111110011101010001111011110111100100000111100011110000110001111011011110100111010010000100111110110100010111100000101101100001000100101001111001111011001101000010010000101011110011000101111101001111011100000000110000011011101001001100010011000110001011110100000011110101010101100110111000111110000010100001011001010000110000110101011111101000111110001001010100100101100001111010101101001011100110101000110101110110000101001101000001011010100000010000101100010010111101111100101000101000110110000001100110100011110011010111011001001000111110101111101100000110011101100000010000111000010010111010001000111100110111010110010111011010111011001010010110010010001101100011010101010011110110101111100111110000000000010000110100001001111101111010010110101001000011110011111011000111011000001001001010111100101010101011100010001100011000101001010110010110001100010101001000100000100011111101000110100110101010110101001100100100000000100111001010101001111111000100000001100111111010000011011010100001001110111011101001111001110000010010000011011110100110100011111110100001000110010101101001101001110010100001011000011101110000010100001110111101110000000101011010111111011110110010110101101001101001110111011110111000110000100111000110101010111000000010110100111000100101100111011100011001101110100001010101111110101000101000000111100100011011000000011101111000001010011101000000101000000010100100011011010101111000001101100011000110101000000000101111110101101001111010101101011000010010110001010000010111100101100111101101101110000010110001111110110001011111010111011000011110000001001110110111010001000001010010110110111110010110101010010111110000110100001110111010110100101111010100110111001110110110010101000001100011101101101110100110110001001101000111101101101001101011111101101010110101000100110000001110111000100000110101010001101010001011010001100110110100010101011000111111001010111001100000100001011000011011110001100111110101011110011011101001100111001100110100000110101111101011001000110001001011001001100110100001101001010001100110001111110110010111101110000010001001111110001010100111110100100101110110110101011010100110010011011011101101010000001001101001001101010110100001101101111101001010001001100100110000010011110010001010011110100001000000010100001100001100101010010111101111011011111001011000011000101001111011100001101010101000010100000111100000110010110111111100100110001011110101100110000000101101101101000110001001101010111001001101010111011010110111101110100011101110011001001000111010100101001110001010011110011010010011101001010101011110011011011000000100001001010111111010111000111100110100110011001110001011111001100110101101111100100110011100111110011110000010100000111011001110011010010101010111100111000010110101000011010010010101110011001101100010111100011100101001110011100110110111001011001111110011001101000010011011001100011110111011001010001100110110101010011011001100011110111100001110111101010111011110010000110100011000110111011101000000010111011110101011000010011111110111010101111000110101001101111010101001111001101011000110001000001001010011000000010111111011011000011001110100011101100000011101111111110010011001000101001101110011001000101101101011111101011111110101100001101001010100101000000110100111010010000001011101101110111101111100001010110011000000110111110001011011100110000011101101011110010010000000101011111100100111110110011111111000101010111110101100001001001011111011011000111001101100000001000101110000001011100101110011110110000011011001101010101101101011111111001011100011001010100111001101111110001011000001110010010110010000001101111111001110100100110100010011100101110111001110110010101010111100011100000110011000110010101000001010110100001001101101100001011011001111010100001001001011111011111001111110101011101010010111000100010101100011001110010111000011010011011100011101100010100000110011110101101110100010111101100110111111101010110110010110110000111111011001111111100000000011100101000010010001000111000101111111000110010000010011000111010000011000110101110010001010110110111111111100001010111010100010111001000111111111110001110100111001000001010001110010000111011110111110001111010000101101011000011110010000111001000011001000110111101110100000110101100010100101000101011100100011010001011000001011110010010000001000110011110010110011110110101101010111100111010111111001000111100111011011101110100111011011011010100110110100010011111010010100000011011000101001100011100100101100010010100111101110010000001001000101110011011010011110110010011011011010111001110111000100010100101000001100110000001101010001011001010110010011100001011010111011010011101110100011110000010110010101011101110000101010101111110010001101101001100001000101101000001111000111000111101011100111101010100100001100111100110111010101010001101010001000010001001111111011011101001000010011111011010111010011000100010001011001100110111100000011111000111010010011000100100111011101000011001000010110000011111100011111001010111101010011101001001000100101100001111101001011111100011010110100100011000010111111111001111101000011110110000011101000100011001100110111010110001111111011001010010101011100001110100101011000011001111000010110110100000001000101101010111111100111010001101100011010011000000011110011101101011001100110110011110010000001011011011000000000110110010001010000100011011110100101110111101111101001100000111100110101000011110111000000011000011101101011011100000100110110100000000100001000110001111101011000110011110101001111110010010001010011010010011101001001111100100010010101110100001010010111011110011010111000111101100011010001011010010100001101101001110110101111001011011101101110110100011010101111010000101010101110110100101000100101111001111110010101110010000111001000001010001001110101000101111100100100101010101101100000000001101111101001011001010101100011111111101010000010011001111100101101110100101001100011110110101111000110100010110001111101000101111000111000001100000110110010011010100011111010111011101011111101110011011111000010001000101000001100000000110000100001010111000100110111110110101000000011001000111101010101000100101101101101010000101010110100111010110101101100111100111111111011111110110011001010110011110000001001011000100110100010011001001001000000100001001100100010000011010111010010001111100001000100101000101001010100100011000111010011111010100110100001011011001010110110001100101101011001100111000011101000111100100111010000111001111110011000101100101001101110100010011000100100001010101011010100010010100101011110000110000000100011101111001001110101110001000100110110110011100110011001000011110110010011001100111010111000010011110110001001001110111010000100000100001000111001000101111100101111000001011001000001010010000111011011000110101001001011000101000111001010101000011111011100111101000010101110100100101000110000001011011000111011010101010001011101010110111001110111010010100100000110011011100101110011100010111011100000101011100110011010010110110101011010000010110011011010001111011111000100110010000011100001001010110000100100100011101000110010000100010001010101011011011110001100001000010000101111010011111101011010000000111110010111101100010100101011011111010100011101110100011011001010010010011011001011011110010101101000000111100010100100101010010100110010110100110100110110111100011111011000010110110001011111000111100110101110000001111000000001001000111010001011110000100001110101111110000101001110111001010001101000000001011001011011100011000111100100010110100010010011000010100100001001001010001111101100100110011100001101001110000110101110000001001010000101110011000111100111111111110101010000010010100111111101101111011110000010000101000111010100111100011100111001100111011111010100000001110001000101001101101010111110101101000011001000010100010110001110101010010110010100000011110111100111111110010000000111001011101000011100010110000101010000000111001111111101101100110001011101011100111010111110011101111110110001101101001011011111010001110011101101000100011000110010110111111101011110110100011010011011011011100111110110110100010000000101000101110110001110011110011101101111110111110011011001100111111111111111010110010111001010101111001110111111110010000001110001000001000111101011011011101100110010111111111000000011000100011011111100010001100111011100111001011001110000000110000111110000110110010011001011101011010000101110110111100110101111111110111101101010000011111101011110111111000011000111001001011100110110000011100001101000000100010100100000011111011110110000110100100100101100011111010000001000111101000100011101001100101011101110110101110011110110111110110110010111111010111001111101011101001110101001000101001110000111001000001100100000110100001111000110010011011001001001011111001110001100000011001001000001001101011100110101011111001001110110111110100011001100001011000000010000110001111110000011101100000100011100100010011110010111111011101100111110100011100100100010011100010011101101010000000100111011001101110001111110110001011011010000110100011100101001110100111001010000000010010101000011110101001110101010000100010110110111011000110010100000001111011010001100001000101110000111101100110010101100000001001001010110001000100001111110110011001101101011011100110001101011100110011001000011100000011000110110001001011010110111111110011000110101111111110000111010010110101111011000011111011000110000111001101110011101100111111100010010011000100100111110100011110001011101010110011111010111111011010011100100011110111101101011101000100110011001010101110001100000100100001111001000011101010011100000101111001011000010011101100110100110011000011100011110110100010110000000001100010100101011000010101111001101010001111000000010110010111101101000011100101110100110000110110100001011000100111010100111111000110100001011111100000110101111011000011110000111111011101101101001110111110010100100000101010100000000110010101110110010011101100110110110000001010110111111110011001111111101101000000010001000010110011000000010101111100001110011000000010010101000100111000100100100111001011100001110100001100111011010101000001011010001010100001101101111110100111100100111100110001110001001110110101110001101111101100000110010011000110011011101100111100101110101101100111001101101101000010010111100111000000011010010111010101101100100100100101111010001111011010010110010011111101000110101110001100010100100010110011001001110001100001010011110010001010010011101111111010011001100011011000101000111111011011000010011101100110000000110010000110001100110100000110011011001010101010110110011100100001000000111101000110010000001000001110101101001111011111000010110110000100011000110111111000101000011101001011110001100001110001111011100010000101001011000011100000100011100000101111001101101110001110110010100110001011100111001011111000001110100000011110001000010000001100010001001011011010000101011001000100101001110101100010010001100000100001110110010111100100110010111111001001001110010101111011000101110101110111110111000011011110110000111001001000111111100000100001110011010000011010010000010001101001000110100010011111010100110001000001110000001000101110111111101111001111110001011110101001111011111100001110100011101000010011110000001000000001101110110111001000111000011000111110000001001101001100011110011011110100111110110000000100010111010101000101000010010001011001010011011000100110111111001100010011101000000000001111110111000110111010011111010010011011010011001101100000111001001100011101111100011110100101001111101100011000100010011111100001001001010010000111111011010111101011011111000110001110001100100001011000000001110101000010100011111110001110100000110100110000010111100010001101100010001100111101010000111100000010011001011110001000000111111111000011000000101111001101000001111100101100101101101110010110001001011010110001100101101111101100001100111111000001100100110111101000101111011001111011100010111010011011010101100110110011000001011000011100010011010101111100110001110111101001110111111001110001011000011011011111100000000001010101100110111101100101000000101001001000000101101101010111000010101010100110011001001111010010001111111100010101111001001111011100000001101110000011101011100011010100001011001110110001010010101100101000010001111111000111010101011001011000000110110011010010101000010111101100011011001001100011000000101000101110101001100110010110100111000001011010110010011001000010100111010000100111011100110111011111000111001010101000001111110110001011110111010101000001110000010010101101100111010000000100011001011000101111100100001010111101011100110101111100011001011010111011111011000000000001100001110110011110110011111010010010010010101101111011000111000011010000100110000010100110000101000111100011111100101100101110011011000001111100111111100111110000110110101100100011001001110011111111101100010010010111000110100010000110010001101011111100110100011110110111101101011110000101010010011001010010011110011111000011100000011001110100001000010000000001111100110100011000110110110100101000000000101111101100010110100010111001001101011011101100100000011100111000101101000110100010111011110110001100111000110000011001010011000111000001100000101111010111010010100001100011111101001111111100101010111111011111000110000101010011110110111000100011011000000000101000000111100000111010110010010110101001001111101000101111101011110001010011111010111011110010101110010001011101010011010001001001100100011100001001000110010010110101111000111100100100111001111100011010100011000011011011001101001101001101111110110110001011000101010101111100000000101100101100001111100101100111011100110001010011111011000101000101110111000101110001111011001000111111110000000100011010100100101111110010000111101110100011100110000000001001100110001101111010000111100111000101000010010101101000110011110100001010011011100001101100111010001001000111100101011001011000011101101100001001100100100101101011010000110101101010101011011010110000010011101100001010100000100100011110001010010000011110001101111101100100101001110111000101001011101101011100010110101011111101110100001100101111100101000101110111011010010001101011110001101000011111001111101000011011110011000101101000000011100110000010010110000001011010100100101111000110111111011010010010000010010001011101000010011001100011011101000000000010000100111111101010101111111010111100010100010000001110101101000100000100000001111011001111110001110001001011100001001111111011101100010110100101101010010001101101001100000111000101100101001011110110010101100011011010001100011000011010100101100100011011001001000101011001010011111000011010100010101000111100111110011011100101101110101110100110101011100101011011101011101100000010011010001111011001111001101010100011101110000000011010001001100011111011011000001010011000110001010010100010001011111001110000001101111001101000001110100101110101110000111001000000111011100110000111110100101110100111111000010101011011000101100101101110011000011101010100101101110110010010001101010101110000010101000001111101011001101111001011110011101101011001000111010110011110110110110110110110001101000110111001001100001001111101110011000101001010010001001011000111101001010000100110010111100010100100000000011000100010100110001110111100011011100110010101001111101011011000110001011111111110110110010110011110101111110100110101111000100001011111111000101000101110100101110010001000100101111110010100101101011001100111110111011001101110001010111011101001101010111001011000001000010100111111101101110001110010010111000000011111011100011100100"
    );

    function h3_get_type(h3type: string; key_width: natural; hash_width: natural) return h3_config;

end package;

package body h3_pack is
    function h3_get_type(h3type: string; key_width: natural; hash_width: natural) return h3_config is
    begin
        if h3type = "AUTO" then
            if key_width <=  H3C_22x11.key_width and hash_width <= H3C_22x11.hash_width then
                return H3C_22x11;
            end if;

            if key_width <=  H3C_64x16.key_width and hash_width <= H3C_64x16.hash_width then
                return H3C_64x16;
            end if;

            if key_width <=  H3C_64x22.key_width and hash_width <= H3C_64x22.hash_width then
                return H3C_64x22;
            end if;

            if key_width <=  H3C_256x64.key_width and hash_width <= H3C_256x64.hash_width then
                return H3C_256x64;
            end if;

            assert false
                report "H3HASH: No hash function was found for given in/out widths! Generate new one using h3_evo tool."
                severity failure;
        else
            if h3type = H3C_22x11.tag then
                return H3C_22x11;
            end if;

            if h3type = H3C_64x16.tag then
                return H3C_64x16;
            end if;

            if h3type = H3C_64x22.tag then
                return H3C_64x22;
            end if;

            if h3type = H3C_256x64.tag then
                return H3C_256x64;
            end if;

            assert false
                report "H3HASH: No hash function was found with the given name!"
                severity failure;
        end if;
    end function;
end package body;

-- watchdog_framelink_ent.vhd: watchdog FrameLink entity
-- Copyright (C) 2015 CESNET
-- Author(s): Adam Piecek <xpiece00@stud.fit.vutbr.cz>
--
-- SPDX-License-Identifier: BSD-3-Clause
--
-- $Id$
--
-- TODO:
--

library IEEE;
use IEEE.std_logic_1164.all;
use WORK.math_pack.all;

entity WATCHDOG_FRAMELINK is
   generic(
      --!   width of the the data flow
      DATA_WIDTH        : positive  := 32;
      --!   enable edge detection on signal KEEP_ALIVE
      EDGE_DETECT       : boolean   := false;
      --!   maximum value of steps to the counter
      COUNT             : positive  := 8;
      --!   width of the counter
      COUNTER_WIDTH     : positive  := 32;
      --!   if TIMING is true, counter counts clock's periods, not data flowing
      TIMING            : boolean   := false
   );

   port(
   -----------------------------------------
   ---        watchdog signals           ---
   -----------------------------------------
      CLK               : in std_logic;
      RESET             : in std_logic;

      --!   counter keep counting
      KEEP_ALIVE        : in std_logic;
      --!   contains exact status of internal counter
      COUNTER           : out std_logic_vector(COUNTER_WIDTH-1 downto 0);
      --!   if watchdog releases data or if it is locked
      LOCKED            : out std_logic;

      -----------------------------------------
      ---        FrameLink signals          ---
      -----------------------------------------

      --! input interface
      RX_DATA             : in  std_logic_vector(DATA_WIDTH-1 downto 0);
      RX_REM              : in  std_logic_vector(LOG2(DATA_WIDTH/8)-1 downto 0);
      RX_SOF_N            : in  std_logic;
      RX_EOF_N            : in  std_logic;
      RX_SOP_N            : in  std_logic;
      RX_EOP_N            : in  std_logic;
      RX_SRC_RDY_IN       : in  std_logic;
      RX_DST_RDY_IN       : out std_logic;

      --! output interface
      TX_DATA             : out std_logic_vector(DATA_WIDTH-1 downto 0);
      TX_REM              : out std_logic_vector(LOG2(DATA_WIDTH/8)-1 downto 0);
      TX_SOF_N            : out std_logic;
      TX_EOF_N            : out std_logic;
      TX_SOP_N            : out std_logic;
      TX_EOP_N            : out std_logic;
      TX_SRC_RDY_OUT      : out std_logic;
      TX_DST_RDY_OUT      : in  std_logic
   );
end;

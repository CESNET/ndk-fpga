//-- data_reg.sv: AVST data register
//-- Copyright (C) 2023 CESNET z. s. p. o.
//-- Author(s): Daniel Kriz <danielkriz@cesnet.cz>

//-- SPDX-License-Identifier: BSD-3-Clause

class data_reg;
    int latency_cnt = 0;
endclass

-- dtb_pack.vhd: DTB Package
-- Copyright (C) 2023 CESNET z. s. p. o.
-- Author(s): Daniel Kriz <danielkriz@cesnet.cz>

-- SPDX-License-Identifier: BSD-3-Clause

library IEEE;
use IEEE.std_logic_1164.all;

package dtb_pkg is

    constant DTB_PF0_DATA : std_logic_vector(8*1272-1 downto 0) := X"5a590100000000028b0d303ee0198876000041f009d10100682865f8000000000000a0d9c2fe81aa42a013e1d9c37eb956e9ea5dd57cef358c782201e48e2f940d00ce01a0ce7374578c9b4cf590c17ab819e12335fa4ab51c0946cc0ace2a2a189d4592ff3b9c4ee6393d5232adadc8804824661e9b65d21036e1b2d8dd430bda67e53872b10f19c53ee98eb34cd799fa27ba6d12346d7b75552aa54bee21344cb94630e49d3af3f76f6b0617bde1a1c9353aafbc43a4774dc20bf1b8e3ed345b1101d52a6069e3b3fbe167479b035a4d195216c7517dd1d0100e8f45ee87bbb0faafe196181ae687f43d1566621c21368e9be3383fd761ef271d2b2d69596de56cf97f4876f7e29b981ac56c1b2ce66573c388ee18f526752254dc205053d96045ef07ae8c4657dc281d636debd90c11e52b42755ac6813453e1d3c09a911168ad2ce8a084e410585b36e2a5e85fa0d6fca9fa261f69d0ead07c80e87be47af834a892dbaf6cf9cfbfe8be9db83156ee81af44e10e4dd22491f5b0d5aecee6539ab1f4fa3949dcede4671dea78f02e11ef700f67e3337f8f87a1cc0820227b01328d73c827ab2c48495f066e46f96831f891732343da60d7c5613b9a4ec09b2e0d6a332e544dc7b2c01fd8bee0e7c891e4e645a3f95a5e3a7acb5ce58959ecbb62bc551274e36b476a9e6f16c675e896b49869ff6d04c4b3b6d8b75b9ee8130d6399da415f4ecf63fc01a46638622124f5437537650339051ab7986c9566be7b523610963854292194d644f23b3def95ff82ca3a95000aa45bea8564009ca31cd8f6c54ee95a85f483588977e209cc41f947c1852240464941335f6dca4855c6cfe793036a15988cdf938c369651486ff926fce5448a33b1478b2bf86c265f72349ac744f78e5e86f62099d506a21691f1424a54dfa1f53417b97a351655b45fda57665833db63f25e3d6d70c29312996d91e9770ad17b663de98c41f1caa21c9dad5b39b88b2d65c23aeb5de271547d24d49b9e145ebcc5213b32979cacf20e1d71d717df6b99433690a0b5a9d0cd9f0f619480ebedef81dd6fd511ec7d4ce42d0ec3e85271553821671114a91a44b0e2611b4b602e5a0b80a0fe3df1dbb9686b0eb91f2a7e1e673f710dec48321f400146cf42035a7ef177d2e842a2395a83a16761ae0e30abc2fbe4a3b98497c5f3a1e124d35cb00fbbc24279bd130ea35f41fa8c4f07c9fd841a3f85080754efb255c0d2da0c8a858a517688635b6317bde92db4c5cb6a218b0b4d5d0a995d6834656a3b35b5716c3e2e5db8bbc4e1a992c48ea3c31ec090e5e8f8e89d854f84ef41c48c37993371d1bb186c5dabd5313bae91533fddc0c564b949c58f578fb6572bf2ad026288fbe767ddbe3d760ce715220d87e5ebd64b015e88231d87c06d15251bcd03576548bc5fff318394f388859f0ff557b496f136242ee98d645ebee8403e2d7f2a1cfef5c7c3634b48a10adee045d96eab352987bc4b2367d1ee141d619065e92b5efbb4969ce2bab4e2bb6bff681768f417dcd6a4e7f16c0afe9c411f44f3a4a9f74b623de40e33bf0f3a705663e565a92e847177af122e25d9e29d882e452448ecca7e6d0eae485635ac40211b272a11712438863bea4087485a0f15b3cec495e2c5594e733b95fadaa7803d030be9d81296deb0bf9a21337220a6bf10d6a2ad14ea8459fef53cddc1fb327ce4c9e57d211c617a25830a8d0f18c95e45d252cd5b0368005db904ef20e0a3e52f74000000160121000236de22690100005a587a37fd";

    constant DTB_VF0_DATA : std_logic_vector(8*0-1 downto 0) := X"";


end package dtb_pkg;

package body dtb_pkg is
end dtb_pkg;
/*
 * sv_flu_pkg.sv: SystemVerilog RMON statistics package
 * Copyright (C) 2016 CESNET
 * Author(s): Pavel Benacek <benacek@cesnet.cz>
 *
 * SPDX-License-Identifier: BSD-3-Clause
 *
 */

package sv_stats_pkg;

  `include "rfc2819_stats.sv"

endpackage : sv_stats_pkg

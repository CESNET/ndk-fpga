/*
 * sv_mi32_pkg.sv: SystemVerilog mi32 package
 * Copyright (C) 2008 CESNET
 * Author(s): Petr Kobiersk� <kobiersky@liberuter.org>
 *            Petr Kastovsky <kastovsky@liberuter.org>
 *
 * SPDX-License-Identifier: BSD-3-Clause
 *
 * $Id$
 *
 * TODO:
 */

// Frame Link Interface
`include "mi32_ifc.sv"

package sv_mi32_pkg;

  import sv_common_pkg::*; // Import SV common classes

  `include "mi32_transaction.sv"
  `include "mi32_driver.sv"
  `include "mi32_monitor.sv"
//  `include "mi32_responder.sv"
//  `include "mi32_command_coverage.sv"

endpackage : sv_mi32_pkg

/*
 * file       : pkg.sv
 * description: test pkg
 * date       : 2020
 * author     : Radek Iša <isa@cesnet.cz>
 *
 * Copyright (C) 2020 CESNET
 * SPDX-License-Identifier: BSD-3-Clause
*/

package test;

    `include "uvm_macros.svh"
    import uvm_pkg::*;

    `include "test.sv"
endpackage
